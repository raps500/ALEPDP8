-- Original: maindec-08-d02b-pb_1-3-68.bin-- This file D02B.vhdl-- CORE memory for the 2100A
--
-- Synchronous read/write block RAM
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity COREMEM is
    port (
        Clock: in  std_logic; 
        ClockEn: in  std_logic; 
        Reset: in  std_logic; 
        WE: in  std_logic; 
        Address: in  std_logic_vector(11 downto 0); 
        Data: in  std_logic_vector(11 downto 0); 
        Q: out  std_logic_vector(11 downto 0)
);

end entity COREMEM;

architecture logic of COREMEM is
    type ram_t is array(natural range 0 to 4095) of std_logic_vector(11 downto 0);
	signal ramdata : ram_t := (
            8#0000# => std_logic_vector(resize(unsigned'(O"5001"), 16)), --             8#0001# => std_logic_vector(resize(unsigned'(O"0002"), 16)), --             8#0002# => std_logic_vector(resize(unsigned'(O"0003"), 16)), --             8#0020# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0021# => std_logic_vector(resize(unsigned'(O"6046"), 16)), --             8#0022# => std_logic_vector(resize(unsigned'(O"6041"), 16)), --             8#0023# => std_logic_vector(resize(unsigned'(O"5022"), 16)), --             8#0024# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#0025# => std_logic_vector(resize(unsigned'(O"5420"), 16)), --             8#0026# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0027# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0030# => std_logic_vector(resize(unsigned'(O"0104"), 16)), --             8#0031# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0032# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0033# => std_logic_vector(resize(unsigned'(O"0103"), 16)), --             8#0034# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0035# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0036# => std_logic_vector(resize(unsigned'(O"0103"), 16)), --             8#0037# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0040# => std_logic_vector(resize(unsigned'(O"5426"), 16)), --             8#0041# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0042# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0043# => std_logic_vector(resize(unsigned'(O"0104"), 16)), --             8#0044# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0045# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0046# => std_logic_vector(resize(unsigned'(O"0103"), 16)), --             8#0047# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0050# => std_logic_vector(resize(unsigned'(O"5441"), 16)), --             8#0051# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0052# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0053# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0054# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0055# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0056# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0057# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0060# => std_logic_vector(resize(unsigned'(O"4000"), 16)), --             8#0061# => std_logic_vector(resize(unsigned'(O"2000"), 16)), --             8#0062# => std_logic_vector(resize(unsigned'(O"1000"), 16)), --             8#0063# => std_logic_vector(resize(unsigned'(O"0400"), 16)), --             8#0064# => std_logic_vector(resize(unsigned'(O"0200"), 16)), --             8#0065# => std_logic_vector(resize(unsigned'(O"0100"), 16)), --             8#0066# => std_logic_vector(resize(unsigned'(O"0040"), 16)), --             8#0067# => std_logic_vector(resize(unsigned'(O"0020"), 16)), --             8#0070# => std_logic_vector(resize(unsigned'(O"0010"), 16)), --             8#0071# => std_logic_vector(resize(unsigned'(O"0004"), 16)), --             8#0072# => std_logic_vector(resize(unsigned'(O"0002"), 16)), --             8#0073# => std_logic_vector(resize(unsigned'(O"0001"), 16)), --             8#0074# => std_logic_vector(resize(unsigned'(O"0057"), 16)), --             8#0075# => std_logic_vector(resize(unsigned'(O"0322"), 16)), --             8#0076# => std_logic_vector(resize(unsigned'(O"0301"), 16)), --             8#0077# => std_logic_vector(resize(unsigned'(O"0314"), 16)), --             8#0100# => std_logic_vector(resize(unsigned'(O"0324"), 16)), --             8#0101# => std_logic_vector(resize(unsigned'(O"0320"), 16)), --             8#0102# => std_logic_vector(resize(unsigned'(O"0240"), 16)), --             8#0103# => std_logic_vector(resize(unsigned'(O"0212"), 16)), --             8#0104# => std_logic_vector(resize(unsigned'(O"0215"), 16)), --             8#0105# => std_logic_vector(resize(unsigned'(O"0060"), 16)), --             8#0106# => std_logic_vector(resize(unsigned'(O"0061"), 16)), --             8#0107# => std_logic_vector(resize(unsigned'(O"0317"), 16)), --             8#0110# => std_logic_vector(resize(unsigned'(O"0313"), 16)), --             8#0111# => std_logic_vector(resize(unsigned'(O"7764"), 16)), --             8#0112# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0113# => std_logic_vector(resize(unsigned'(O"0262"), 16)), --             8#0114# => std_logic_vector(resize(unsigned'(O"0302"), 16)), --             8#0115# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0116# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0117# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0120# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0121# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0122# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0123# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0124# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0125# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0126# => std_logic_vector(resize(unsigned'(O"7776"), 16)), --             8#0127# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0130# => std_logic_vector(resize(unsigned'(O"0307"), 16)), --             8#0131# => std_logic_vector(resize(unsigned'(O"0304"), 16)), --             8#0132# => std_logic_vector(resize(unsigned'(O"0330"), 16)), --             8#0133# => std_logic_vector(resize(unsigned'(O"0331"), 16)), --             8#0134# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0135# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0136# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0137# => std_logic_vector(resize(unsigned'(O"7763"), 16)), --             8#0140# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0141# => std_logic_vector(resize(unsigned'(O"7377"), 16)), --             8#0142# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0143# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0144# => std_logic_vector(resize(unsigned'(O"0140"), 16)), --             8#0145# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0146# => std_logic_vector(resize(unsigned'(O"5150"), 16)), --             8#0147# => std_logic_vector(resize(unsigned'(O"5152"), 16)), --             8#0150# => std_logic_vector(resize(unsigned'(O"7360"), 16)), --             8#0151# => std_logic_vector(resize(unsigned'(O"5542"), 16)), --             8#0152# => std_logic_vector(resize(unsigned'(O"7340"), 16)), --             8#0153# => std_logic_vector(resize(unsigned'(O"5542"), 16)), --             8#0000# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#0001# => std_logic_vector(resize(unsigned'(O"1417"), 16)), --             8#0002# => std_logic_vector(resize(unsigned'(O"3135"), 16)), --             8#0003# => std_logic_vector(resize(unsigned'(O"1417"), 16)), --             8#0004# => std_logic_vector(resize(unsigned'(O"3136"), 16)), --             8#0005# => std_logic_vector(resize(unsigned'(O"2216"), 16)), --             8#0006# => std_logic_vector(resize(unsigned'(O"5647"), 16)), --             8#0007# => std_logic_vector(resize(unsigned'(O"1215"), 16)), --             8#0010# => std_logic_vector(resize(unsigned'(O"3017"), 16)), --             8#0011# => std_logic_vector(resize(unsigned'(O"1214"), 16)), --             8#0012# => std_logic_vector(resize(unsigned'(O"3216"), 16)), --             8#0013# => std_logic_vector(resize(unsigned'(O"5647"), 16)), --             8#0014# => std_logic_vector(resize(unsigned'(O"7634"), 16)), --             8#0015# => std_logic_vector(resize(unsigned'(O"4177"), 16)), --             8#0016# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0017# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0020# => std_logic_vector(resize(unsigned'(O"7300"), 16)), --             8#0021# => std_logic_vector(resize(unsigned'(O"2217"), 16)), --             8#0022# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0023# => std_logic_vector(resize(unsigned'(O"1217"), 16)), --             8#0024# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#0025# => std_logic_vector(resize(unsigned'(O"7630"), 16)), --             8#0026# => std_logic_vector(resize(unsigned'(O"5230"), 16)), --             8#0027# => std_logic_vector(resize(unsigned'(O"5200"), 16)), --             8#0030# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#0031# => std_logic_vector(resize(unsigned'(O"0063"), 16)), --             8#0032# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0033# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0034# => std_logic_vector(resize(unsigned'(O"5650"), 16)), --             8#0035# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0036# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#0037# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0040# => std_logic_vector(resize(unsigned'(O"3135"), 16)), --             8#0041# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0042# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#0043# => std_logic_vector(resize(unsigned'(O"7001"), 16)), --             8#0044# => std_logic_vector(resize(unsigned'(O"1410"), 16)), --             8#0045# => std_logic_vector(resize(unsigned'(O"3136"), 16)), --             8#0046# => std_logic_vector(resize(unsigned'(O"5647"), 16)), --             8#0047# => std_logic_vector(resize(unsigned'(O"0225"), 16)), --             8#0050# => std_logic_vector(resize(unsigned'(O"0312"), 16)), --             8#0017# => std_logic_vector(resize(unsigned'(O"4177"), 16)), --             8#0051# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0052# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#0053# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0054# => std_logic_vector(resize(unsigned'(O"0122"), 16)), --             8#0055# => std_logic_vector(resize(unsigned'(O"3275"), 16)), --             8#0056# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0057# => std_logic_vector(resize(unsigned'(O"0122"), 16)), --             8#0060# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0061# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#0062# => std_logic_vector(resize(unsigned'(O"3274"), 16)), --             8#0063# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0064# => std_logic_vector(resize(unsigned'(O"0275"), 16)), --             8#0065# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0066# => std_logic_vector(resize(unsigned'(O"5676"), 16)), --             8#0067# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0070# => std_logic_vector(resize(unsigned'(O"0274"), 16)), --             8#0071# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0072# => std_logic_vector(resize(unsigned'(O"5676"), 16)), --             8#0073# => std_logic_vector(resize(unsigned'(O"5277"), 16)), --             8#0074# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0075# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0076# => std_logic_vector(resize(unsigned'(O"0400"), 16)), --             8#0077# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0100# => std_logic_vector(resize(unsigned'(O"0134"), 16)), --             8#0101# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0102# => std_logic_vector(resize(unsigned'(O"0120"), 16)), --             8#0103# => std_logic_vector(resize(unsigned'(O"3322"), 16)), --             8#0104# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0105# => std_logic_vector(resize(unsigned'(O"0120"), 16)), --             8#0106# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0107# => std_logic_vector(resize(unsigned'(O"0134"), 16)), --             8#0110# => std_logic_vector(resize(unsigned'(O"3323"), 16)), --             8#0111# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0112# => std_logic_vector(resize(unsigned'(O"0322"), 16)), --             8#0113# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0114# => std_logic_vector(resize(unsigned'(O"5676"), 16)), --             8#0115# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0116# => std_logic_vector(resize(unsigned'(O"0323"), 16)), --             8#0117# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0120# => std_logic_vector(resize(unsigned'(O"5676"), 16)), --             8#0121# => std_logic_vector(resize(unsigned'(O"5724"), 16)), --             8#0122# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0123# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0124# => std_logic_vector(resize(unsigned'(O"0407"), 16)), --             8#1000# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1001# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1002# => std_logic_vector(resize(unsigned'(O"7776"), 16)), --             8#1003# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1004# => std_logic_vector(resize(unsigned'(O"7775"), 16)), --             8#1005# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1006# => std_logic_vector(resize(unsigned'(O"7773"), 16)), --             8#1007# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1010# => std_logic_vector(resize(unsigned'(O"7767"), 16)), --             8#1011# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1012# => std_logic_vector(resize(unsigned'(O"7757"), 16)), --             8#1013# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1014# => std_logic_vector(resize(unsigned'(O"7737"), 16)), --             8#1015# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1016# => std_logic_vector(resize(unsigned'(O"7677"), 16)), --             8#1017# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1020# => std_logic_vector(resize(unsigned'(O"7577"), 16)), --             8#1021# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1022# => std_logic_vector(resize(unsigned'(O"7377"), 16)), --             8#1023# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1024# => std_logic_vector(resize(unsigned'(O"6777"), 16)), --             8#1025# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1026# => std_logic_vector(resize(unsigned'(O"5777"), 16)), --             8#1027# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1030# => std_logic_vector(resize(unsigned'(O"3777"), 16)), --             8#1031# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1032# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1033# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1034# => std_logic_vector(resize(unsigned'(O"7776"), 16)), --             8#1035# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1036# => std_logic_vector(resize(unsigned'(O"7775"), 16)), --             8#1037# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1040# => std_logic_vector(resize(unsigned'(O"7773"), 16)), --             8#1041# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1042# => std_logic_vector(resize(unsigned'(O"7767"), 16)), --             8#1043# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1044# => std_logic_vector(resize(unsigned'(O"7757"), 16)), --             8#1045# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1046# => std_logic_vector(resize(unsigned'(O"7737"), 16)), --             8#1047# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1050# => std_logic_vector(resize(unsigned'(O"7677"), 16)), --             8#1051# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1052# => std_logic_vector(resize(unsigned'(O"7577"), 16)), --             8#1053# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1054# => std_logic_vector(resize(unsigned'(O"7377"), 16)), --             8#1055# => std_logic_vector(resize(unsigned'(O"6777"), 16)), --             8#1056# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1057# => std_logic_vector(resize(unsigned'(O"5777"), 16)), --             8#1060# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1061# => std_logic_vector(resize(unsigned'(O"3777"), 16)), --             8#1062# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1063# => std_logic_vector(resize(unsigned'(O"0001"), 16)), --             8#1064# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1065# => std_logic_vector(resize(unsigned'(O"0002"), 16)), --             8#1066# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1067# => std_logic_vector(resize(unsigned'(O"0004"), 16)), --             8#1070# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1071# => std_logic_vector(resize(unsigned'(O"0010"), 16)), --             8#1072# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1073# => std_logic_vector(resize(unsigned'(O"0020"), 16)), --             8#1074# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1075# => std_logic_vector(resize(unsigned'(O"0040"), 16)), --             8#1076# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1077# => std_logic_vector(resize(unsigned'(O"0100"), 16)), --             8#1100# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1101# => std_logic_vector(resize(unsigned'(O"0200"), 16)), --             8#1102# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1103# => std_logic_vector(resize(unsigned'(O"0400"), 16)), --             8#1104# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1105# => std_logic_vector(resize(unsigned'(O"1000"), 16)), --             8#1106# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1107# => std_logic_vector(resize(unsigned'(O"2000"), 16)), --             8#1110# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1111# => std_logic_vector(resize(unsigned'(O"4000"), 16)), --             8#1112# => std_logic_vector(resize(unsigned'(O"0001"), 16)), --             8#1113# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1114# => std_logic_vector(resize(unsigned'(O"0002"), 16)), --             8#1115# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1116# => std_logic_vector(resize(unsigned'(O"0004"), 16)), --             8#1117# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1120# => std_logic_vector(resize(unsigned'(O"0010"), 16)), --             8#1121# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1122# => std_logic_vector(resize(unsigned'(O"0200"), 16)), --             8#1123# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1124# => std_logic_vector(resize(unsigned'(O"0400"), 16)), --             8#1125# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1126# => std_logic_vector(resize(unsigned'(O"0100"), 16)), --             8#1127# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1130# => std_logic_vector(resize(unsigned'(O"0200"), 16)), --             8#1131# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1132# => std_logic_vector(resize(unsigned'(O"0400"), 16)), --             8#1133# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1134# => std_logic_vector(resize(unsigned'(O"1000"), 16)), --             8#1135# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1136# => std_logic_vector(resize(unsigned'(O"2000"), 16)), --             8#1137# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1140# => std_logic_vector(resize(unsigned'(O"4000"), 16)), --             8#1141# => std_logic_vector(resize(unsigned'(O"7777"), 16)), --             8#1000# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1001# => std_logic_vector(resize(unsigned'(O"3124"), 16)), --             8#1002# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1003# => std_logic_vector(resize(unsigned'(O"3135"), 16)), --             8#1004# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1005# => std_logic_vector(resize(unsigned'(O"3136"), 16)), --             8#1006# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1007# => std_logic_vector(resize(unsigned'(O"3121"), 16)), --             8#1010# => std_logic_vector(resize(unsigned'(O"3134"), 16)), --             8#1011# => std_logic_vector(resize(unsigned'(O"3115"), 16)), --             8#1012# => std_logic_vector(resize(unsigned'(O"5223"), 16)), --             8#1013# => std_logic_vector(resize(unsigned'(O"3120"), 16)), --             8#1014# => std_logic_vector(resize(unsigned'(O"7340"), 16)), --             8#1015# => std_logic_vector(resize(unsigned'(O"0135"), 16)), --             8#1016# => std_logic_vector(resize(unsigned'(O"1136"), 16)), --             8#1017# => std_logic_vector(resize(unsigned'(O"3122"), 16)), --             8#1020# => std_logic_vector(resize(unsigned'(O"7004"), 16)), --             8#1021# => std_logic_vector(resize(unsigned'(O"3134"), 16)), --             8#1022# => std_logic_vector(resize(unsigned'(O"5737"), 16)), --             8#1023# => std_logic_vector(resize(unsigned'(O"5624"), 16)), --             8#1024# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1025# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1026# => std_logic_vector(resize(unsigned'(O"0135"), 16)), --             8#1027# => std_logic_vector(resize(unsigned'(O"3115"), 16)), --             8#1030# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1031# => std_logic_vector(resize(unsigned'(O"0136"), 16)), --             8#1032# => std_logic_vector(resize(unsigned'(O"3116"), 16)), --             8#1033# => std_logic_vector(resize(unsigned'(O"4235"), 16)), --             8#1034# => std_logic_vector(resize(unsigned'(O"5214"), 16)), --             8#1035# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#1036# => std_logic_vector(resize(unsigned'(O"7300"), 16)), --             8#1037# => std_logic_vector(resize(unsigned'(O"3121"), 16)), --             8#1040# => std_logic_vector(resize(unsigned'(O"3120"), 16)), --             8#1041# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1042# => std_logic_vector(resize(unsigned'(O"0111"), 16)), --             8#1043# => std_logic_vector(resize(unsigned'(O"3123"), 16)), --             8#1044# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1045# => std_logic_vector(resize(unsigned'(O"0115"), 16)), --             8#1046# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#1047# => std_logic_vector(resize(unsigned'(O"3115"), 16)), --             8#1050# => std_logic_vector(resize(unsigned'(O"7004"), 16)), --             8#1051# => std_logic_vector(resize(unsigned'(O"3117"), 16)), --             8#1052# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1053# => std_logic_vector(resize(unsigned'(O"0116"), 16)), --             8#1054# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#1055# => std_logic_vector(resize(unsigned'(O"3116"), 16)), --             8#1056# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1057# => std_logic_vector(resize(unsigned'(O"0117"), 16)), --             8#1060# => std_logic_vector(resize(unsigned'(O"7420"), 16)), --             8#1061# => std_logic_vector(resize(unsigned'(O"5302"), 16)), --             8#1062# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#1063# => std_logic_vector(resize(unsigned'(O"5305"), 16)), --             8#1064# => std_logic_vector(resize(unsigned'(O"7300"), 16)), --             8#1065# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1066# => std_logic_vector(resize(unsigned'(O"0120"), 16)), --             8#1067# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#1070# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1071# => std_logic_vector(resize(unsigned'(O"0117"), 16)), --             8#1072# => std_logic_vector(resize(unsigned'(O"3120"), 16)), --             8#1073# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1074# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#1075# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#1076# => std_logic_vector(resize(unsigned'(O"3121"), 16)), --             8#1077# => std_logic_vector(resize(unsigned'(O"2123"), 16)), --             8#1100# => std_logic_vector(resize(unsigned'(O"5244"), 16)), --             8#1101# => std_logic_vector(resize(unsigned'(O"5635"), 16)), --             8#1102# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#1103# => std_logic_vector(resize(unsigned'(O"5265"), 16)), --             8#1104# => std_logic_vector(resize(unsigned'(O"7220"), 16)), --             8#1105# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1106# => std_logic_vector(resize(unsigned'(O"0120"), 16)), --             8#1107# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#1110# => std_logic_vector(resize(unsigned'(O"7100"), 16)), --             8#1111# => std_logic_vector(resize(unsigned'(O"5272"), 16)), --             8#1112# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#1113# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1114# => std_logic_vector(resize(unsigned'(O"0076"), 16)), --             8#1115# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1116# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1117# => std_logic_vector(resize(unsigned'(O"0131"), 16)), --             8#1120# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1121# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1122# => std_logic_vector(resize(unsigned'(O"0131"), 16)), --             8#1123# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1124# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1125# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#1126# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1127# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1130# => std_logic_vector(resize(unsigned'(O"0107"), 16)), --             8#1131# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1132# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#1133# => std_logic_vector(resize(unsigned'(O"0110"), 16)), --             8#1134# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#1135# => std_logic_vector(resize(unsigned'(O"5736"), 16)), --             8#1136# => std_logic_vector(resize(unsigned'(O"2000"), 16)), --             8#1137# => std_logic_vector(resize(unsigned'(O"4051"), 16)), --             8#2000# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2001# => std_logic_vector(resize(unsigned'(O"7106"), 16)), --             8#2002# => std_logic_vector(resize(unsigned'(O"7510"), 16)), --             8#2003# => std_logic_vector(resize(unsigned'(O"4216"), 16)), --             8#2004# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2005# => std_logic_vector(resize(unsigned'(O"7510"), 16)), --             8#2006# => std_logic_vector(resize(unsigned'(O"7402"), 16)), --             8#2007# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2010# => std_logic_vector(resize(unsigned'(O"7104"), 16)), --             8#2011# => std_logic_vector(resize(unsigned'(O"7510"), 16)), --             8#2012# => std_logic_vector(resize(unsigned'(O"5614"), 16)), --             8#2013# => std_logic_vector(resize(unsigned'(O"5615"), 16)), --             8#2014# => std_logic_vector(resize(unsigned'(O"0225"), 16)), --             8#2015# => std_logic_vector(resize(unsigned'(O"0223"), 16)), --             8#2016# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2017# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2020# => std_logic_vector(resize(unsigned'(O"0124"), 16)), --             8#2021# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#2022# => std_logic_vector(resize(unsigned'(O"4321"), 16)), --             8#2023# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#2024# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#2025# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2026# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2027# => std_logic_vector(resize(unsigned'(O"0120"), 16)), --             8#2030# => std_logic_vector(resize(unsigned'(O"4635"), 16)), --             8#2031# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2032# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#2033# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2034# => std_logic_vector(resize(unsigned'(O"5236"), 16)), --             8#2035# => std_logic_vector(resize(unsigned'(O"2637"), 16)), --             8#2036# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2037# => std_logic_vector(resize(unsigned'(O"0121"), 16)), --             8#2040# => std_logic_vector(resize(unsigned'(O"3125"), 16)), --             8#2041# => std_logic_vector(resize(unsigned'(O"4266"), 16)), --             8#2042# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2043# => std_logic_vector(resize(unsigned'(O"0134"), 16)), --             8#2044# => std_logic_vector(resize(unsigned'(O"4635"), 16)), --             8#2045# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2046# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#2047# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2050# => std_logic_vector(resize(unsigned'(O"5251"), 16)), --             8#2051# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2052# => std_logic_vector(resize(unsigned'(O"0122"), 16)), --             8#2053# => std_logic_vector(resize(unsigned'(O"3125"), 16)), --             8#2054# => std_logic_vector(resize(unsigned'(O"4266"), 16)), --             8#2055# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2056# => std_logic_vector(resize(unsigned'(O"0135"), 16)), --             8#2057# => std_logic_vector(resize(unsigned'(O"3125"), 16)), --             8#2060# => std_logic_vector(resize(unsigned'(O"4266"), 16)), --             8#2061# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2062# => std_logic_vector(resize(unsigned'(O"0136"), 16)), --             8#2063# => std_logic_vector(resize(unsigned'(O"3125"), 16)), --             8#2064# => std_logic_vector(resize(unsigned'(O"4266"), 16)), --             8#2065# => std_logic_vector(resize(unsigned'(O"5616"), 16)), --             8#2066# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2067# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2070# => std_logic_vector(resize(unsigned'(O"0137"), 16)), --             8#2071# => std_logic_vector(resize(unsigned'(O"3112"), 16)), --             8#2072# => std_logic_vector(resize(unsigned'(O"2112"), 16)), --             8#2073# => std_logic_vector(resize(unsigned'(O"7410"), 16)), --             8#2074# => std_logic_vector(resize(unsigned'(O"5312"), 16)), --             8#2075# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2076# => std_logic_vector(resize(unsigned'(O"0125"), 16)), --             8#2077# => std_logic_vector(resize(unsigned'(O"7100"), 16)), --             8#2100# => std_logic_vector(resize(unsigned'(O"7004"), 16)), --             8#2101# => std_logic_vector(resize(unsigned'(O"3125"), 16)), --             8#2102# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#2103# => std_logic_vector(resize(unsigned'(O"5306"), 16)), --             8#2104# => std_logic_vector(resize(unsigned'(O"4764"), 16)), --             8#2105# => std_logic_vector(resize(unsigned'(O"5272"), 16)), --             8#2106# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2107# => std_logic_vector(resize(unsigned'(O"0106"), 16)), --             8#2110# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2111# => std_logic_vector(resize(unsigned'(O"5272"), 16)), --             8#2112# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2113# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#2114# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2115# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2116# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#2117# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2120# => std_logic_vector(resize(unsigned'(O"5666"), 16)), --             8#2121# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2122# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2123# => std_logic_vector(resize(unsigned'(O"3124"), 16)), --             8#2124# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2125# => std_logic_vector(resize(unsigned'(O"0126"), 16)), --             8#2126# => std_logic_vector(resize(unsigned'(O"3127"), 16)), --             8#2127# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#2130# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2131# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#2132# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2133# => std_logic_vector(resize(unsigned'(O"2127"), 16)), --             8#2134# => std_logic_vector(resize(unsigned'(O"5330"), 16)), --             8#2135# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2136# => std_logic_vector(resize(unsigned'(O"0130"), 16)), --             8#2137# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2140# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2141# => std_logic_vector(resize(unsigned'(O"0107"), 16)), --             8#2142# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2143# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2144# => std_logic_vector(resize(unsigned'(O"0107"), 16)), --             8#2145# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2146# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2147# => std_logic_vector(resize(unsigned'(O"0131"), 16)), --             8#2150# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2151# => std_logic_vector(resize(unsigned'(O"4762"), 16)), --             8#2152# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2153# => std_logic_vector(resize(unsigned'(O"0114"), 16)), --             8#2154# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2155# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#2156# => std_logic_vector(resize(unsigned'(O"0076"), 16)), --             8#2157# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2160# => std_logic_vector(resize(unsigned'(O"5761"), 16)), --             8#2161# => std_logic_vector(resize(unsigned'(O"0600"), 16)), --             8#2162# => std_logic_vector(resize(unsigned'(O"0626"), 16)), --             8#2163# => std_logic_vector(resize(unsigned'(O"5721"), 16)), --             8#2164# => std_logic_vector(resize(unsigned'(O"2702"), 16)), --             8#3000# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3001# => std_logic_vector(resize(unsigned'(O"0131"), 16)), --             8#3002# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3003# => std_logic_vector(resize(unsigned'(O"4226"), 16)), --             8#3004# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3005# => std_logic_vector(resize(unsigned'(O"0132"), 16)), --             8#3006# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3007# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3010# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#3011# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3012# => std_logic_vector(resize(unsigned'(O"4240"), 16)), --             8#3013# => std_logic_vector(resize(unsigned'(O"4226"), 16)), --             8#3014# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3015# => std_logic_vector(resize(unsigned'(O"0133"), 16)), --             8#3016# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3017# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3020# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#3021# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3022# => std_logic_vector(resize(unsigned'(O"4240"), 16)), --             8#3023# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#3024# => std_logic_vector(resize(unsigned'(O"5625"), 16)), --             8#3025# => std_logic_vector(resize(unsigned'(O"0563"), 16)), --             8#3026# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3027# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3030# => std_logic_vector(resize(unsigned'(O"0111"), 16)), --             8#3031# => std_logic_vector(resize(unsigned'(O"3127"), 16)), --             8#3032# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3033# => std_logic_vector(resize(unsigned'(O"0102"), 16)), --             8#3034# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3035# => std_logic_vector(resize(unsigned'(O"2127"), 16)), --             8#3036# => std_logic_vector(resize(unsigned'(O"5232"), 16)), --             8#3037# => std_logic_vector(resize(unsigned'(O"5626"), 16)), --             8#3040# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3041# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3042# => std_logic_vector(resize(unsigned'(O"0076"), 16)), --             8#3043# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3044# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3045# => std_logic_vector(resize(unsigned'(O"0075"), 16)), --             8#3046# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3047# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3050# => std_logic_vector(resize(unsigned'(O"0130"), 16)), --             8#3051# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3052# => std_logic_vector(resize(unsigned'(O"5640"), 16)), --             8#0000# => std_logic_vector(resize(unsigned'(O"4316"), 16)), --             8#0001# => std_logic_vector(resize(unsigned'(O"4142"), 16)), --             8#0002# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0003# => std_logic_vector(resize(unsigned'(O"7001"), 16)), --             8#0004# => std_logic_vector(resize(unsigned'(O"3051"), 16)), --             8#0005# => std_logic_vector(resize(unsigned'(O"7420"), 16)), --             8#0006# => std_logic_vector(resize(unsigned'(O"5215"), 16)), --             8#0007# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#0010# => std_logic_vector(resize(unsigned'(O"3140"), 16)), --             8#0011# => std_logic_vector(resize(unsigned'(O"4352"), 16)), --             8#0012# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0013# => std_logic_vector(resize(unsigned'(O"5220"), 16)), --             8#0014# => std_logic_vector(resize(unsigned'(O"5274"), 16)), --             8#0015# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#0016# => std_logic_vector(resize(unsigned'(O"3140"), 16)), --             8#0017# => std_logic_vector(resize(unsigned'(O"5211"), 16)), --             8#0020# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0021# => std_logic_vector(resize(unsigned'(O"3056"), 16)), --             8#0022# => std_logic_vector(resize(unsigned'(O"7340"), 16)), --             8#0023# => std_logic_vector(resize(unsigned'(O"0140"), 16)), --             8#0024# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0025# => std_logic_vector(resize(unsigned'(O"5272"), 16)), --             8#0026# => std_logic_vector(resize(unsigned'(O"7140"), 16)), --             8#0027# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0030# => std_logic_vector(resize(unsigned'(O"7004"), 16)), --             8#0031# => std_logic_vector(resize(unsigned'(O"3052"), 16)), --             8#0032# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#0033# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#0034# => std_logic_vector(resize(unsigned'(O"3053"), 16)), --             8#0035# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0036# => std_logic_vector(resize(unsigned'(O"0052"), 16)), --             8#0037# => std_logic_vector(resize(unsigned'(O"7010"), 16)), --             8#0040# => std_logic_vector(resize(unsigned'(O"3054"), 16)), --             8#0041# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#0042# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#0043# => std_logic_vector(resize(unsigned'(O"3055"), 16)), --             8#0044# => std_logic_vector(resize(unsigned'(O"7340"), 16)), --             8#0045# => std_logic_vector(resize(unsigned'(O"0054"), 16)), --             8#0046# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0047# => std_logic_vector(resize(unsigned'(O"1051"), 16)), --             8#0050# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0051# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#0052# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#0053# => std_logic_vector(resize(unsigned'(O"5715"), 16)), --             8#0054# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#0055# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0056# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0057# => std_logic_vector(resize(unsigned'(O"1053"), 16)), --             8#0060# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0061# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0062# => std_logic_vector(resize(unsigned'(O"5715"), 16)), --             8#0063# => std_logic_vector(resize(unsigned'(O"1055"), 16)), --             8#0064# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0065# => std_logic_vector(resize(unsigned'(O"1140"), 16)), --             8#0066# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0067# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0070# => std_logic_vector(resize(unsigned'(O"5715"), 16)), --             8#0071# => std_logic_vector(resize(unsigned'(O"5751"), 16)), --             8#0072# => std_logic_vector(resize(unsigned'(O"7360"), 16)), --             8#0073# => std_logic_vector(resize(unsigned'(O"5227"), 16)), --             8#0074# => std_logic_vector(resize(unsigned'(O"4316"), 16)), --             8#0075# => std_logic_vector(resize(unsigned'(O"4142"), 16)), --             8#0076# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0077# => std_logic_vector(resize(unsigned'(O"7001"), 16)), --             8#0100# => std_logic_vector(resize(unsigned'(O"3051"), 16)), --             8#0101# => std_logic_vector(resize(unsigned'(O"7420"), 16)), --             8#0102# => std_logic_vector(resize(unsigned'(O"5311"), 16)), --             8#0103# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#0104# => std_logic_vector(resize(unsigned'(O"3140"), 16)), --             8#0105# => std_logic_vector(resize(unsigned'(O"4363"), 16)), --             8#0106# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0107# => std_logic_vector(resize(unsigned'(O"5714"), 16)), --             8#0110# => std_logic_vector(resize(unsigned'(O"5332"), 16)), --             8#0111# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#0112# => std_logic_vector(resize(unsigned'(O"3140"), 16)), --             8#0113# => std_logic_vector(resize(unsigned'(O"5305"), 16)), --             8#0114# => std_logic_vector(resize(unsigned'(O"2200"), 16)), --             8#0115# => std_logic_vector(resize(unsigned'(O"2400"), 16)), --             8#0116# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0117# => std_logic_vector(resize(unsigned'(O"7300"), 16)), --             8#0120# => std_logic_vector(resize(unsigned'(O"3051"), 16)), --             8#0121# => std_logic_vector(resize(unsigned'(O"3052"), 16)), --             8#0122# => std_logic_vector(resize(unsigned'(O"3054"), 16)), --             8#0123# => std_logic_vector(resize(unsigned'(O"3053"), 16)), --             8#0124# => std_logic_vector(resize(unsigned'(O"3055"), 16)), --             8#0125# => std_logic_vector(resize(unsigned'(O"3140"), 16)), --             8#0126# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0127# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0130# => std_logic_vector(resize(unsigned'(O"7000"), 16)), --             8#0131# => std_logic_vector(resize(unsigned'(O"5716"), 16)), --             8#0132# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#0133# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#0134# => std_logic_vector(resize(unsigned'(O"1075"), 16)), --             8#0135# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0136# => std_logic_vector(resize(unsigned'(O"1107"), 16)), --             8#0137# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0140# => std_logic_vector(resize(unsigned'(O"1100"), 16)), --             8#0141# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0142# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#0143# => std_logic_vector(resize(unsigned'(O"1113"), 16)), --             8#0144# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0145# => std_logic_vector(resize(unsigned'(O"1114"), 16)), --             8#0146# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#0147# => std_logic_vector(resize(unsigned'(O"5750"), 16)), --             8#0150# => std_logic_vector(resize(unsigned'(O"0200"), 16)), --             8#0151# => std_logic_vector(resize(unsigned'(O"2521"), 16)), --             8#0152# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0153# => std_logic_vector(resize(unsigned'(O"1140"), 16)), --             8#0154# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0155# => std_logic_vector(resize(unsigned'(O"7410"), 16)), --             8#0156# => std_logic_vector(resize(unsigned'(O"5220"), 16)), --             8#0157# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0160# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0161# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0162# => std_logic_vector(resize(unsigned'(O"5752"), 16)), --             8#0163# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0164# => std_logic_vector(resize(unsigned'(O"1140"), 16)), --             8#0165# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#0166# => std_logic_vector(resize(unsigned'(O"7410"), 16)), --             8#0167# => std_logic_vector(resize(unsigned'(O"5714"), 16)), --             8#0170# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#0171# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#0172# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#0173# => std_logic_vector(resize(unsigned'(O"5763"), 16)), --             8#1000# => std_logic_vector(resize(unsigned'(O"7300"), 16)), --             8#1001# => std_logic_vector(resize(unsigned'(O"3056"), 16)), --             8#1002# => std_logic_vector(resize(unsigned'(O"7340"), 16)), --             8#1003# => std_logic_vector(resize(unsigned'(O"0140"), 16)), --             8#1004# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#1005# => std_logic_vector(resize(unsigned'(O"5250"), 16)), --             8#1006# => std_logic_vector(resize(unsigned'(O"7140"), 16)), --             8#1007# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#1010# => std_logic_vector(resize(unsigned'(O"7012"), 16)), --             8#1011# => std_logic_vector(resize(unsigned'(O"3054"), 16)), --             8#1012# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#1013# => std_logic_vector(resize(unsigned'(O"1072"), 16)), --             8#1014# => std_logic_vector(resize(unsigned'(O"3055"), 16)), --             8#1015# => std_logic_vector(resize(unsigned'(O"1054"), 16)), --             8#1016# => std_logic_vector(resize(unsigned'(O"7006"), 16)), --             8#1017# => std_logic_vector(resize(unsigned'(O"3052"), 16)), --             8#1020# => std_logic_vector(resize(unsigned'(O"7430"), 16)), --             8#1021# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#1022# => std_logic_vector(resize(unsigned'(O"3053"), 16)), --             8#1023# => std_logic_vector(resize(unsigned'(O"7100"), 16)), --             8#1024# => std_logic_vector(resize(unsigned'(O"1052"), 16)), --             8#1025# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1026# => std_logic_vector(resize(unsigned'(O"1051"), 16)), --             8#1027# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1030# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#1031# => std_logic_vector(resize(unsigned'(O"5652"), 16)), --             8#1032# => std_logic_vector(resize(unsigned'(O"1072"), 16)), --             8#1033# => std_logic_vector(resize(unsigned'(O"0051"), 16)), --             8#1034# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1035# => std_logic_vector(resize(unsigned'(O"1055"), 16)), --             8#1036# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1037# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#1040# => std_logic_vector(resize(unsigned'(O"5652"), 16)), --             8#1041# => std_logic_vector(resize(unsigned'(O"1053"), 16)), --             8#1042# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1043# => std_logic_vector(resize(unsigned'(O"1140"), 16)), --             8#1044# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#1045# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#1046# => std_logic_vector(resize(unsigned'(O"5652"), 16)), --             8#1047# => std_logic_vector(resize(unsigned'(O"5653"), 16)), --             8#1050# => std_logic_vector(resize(unsigned'(O"7360"), 16)), --             8#1051# => std_logic_vector(resize(unsigned'(O"5207"), 16)), --             8#1052# => std_logic_vector(resize(unsigned'(O"2406"), 16)), --             8#1053# => std_logic_vector(resize(unsigned'(O"2525"), 16)), --             8#2000# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2001# => std_logic_vector(resize(unsigned'(O"1244"), 16)), --             8#2002# => std_logic_vector(resize(unsigned'(O"3215"), 16)), --             8#2003# => std_logic_vector(resize(unsigned'(O"1245"), 16)), --             8#2004# => std_logic_vector(resize(unsigned'(O"3214"), 16)), --             8#2005# => std_logic_vector(resize(unsigned'(O"5216"), 16)), --             8#2006# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2007# => std_logic_vector(resize(unsigned'(O"1250"), 16)), --             8#2010# => std_logic_vector(resize(unsigned'(O"3215"), 16)), --             8#2011# => std_logic_vector(resize(unsigned'(O"1251"), 16)), --             8#2012# => std_logic_vector(resize(unsigned'(O"3214"), 16)), --             8#2013# => std_logic_vector(resize(unsigned'(O"5216"), 16)), --             8#2014# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2015# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2016# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2017# => std_logic_vector(resize(unsigned'(O"0062"), 16)), --             8#2020# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2021# => std_logic_vector(resize(unsigned'(O"1062"), 16)), --             8#2022# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2023# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#2024# => std_logic_vector(resize(unsigned'(O"4255"), 16)), --             8#2025# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2026# => std_logic_vector(resize(unsigned'(O"0060"), 16)), --             8#2027# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2030# => std_logic_vector(resize(unsigned'(O"1060"), 16)), --             8#2031# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2032# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#2033# => std_logic_vector(resize(unsigned'(O"7402"), 16)), --             8#2034# => std_logic_vector(resize(unsigned'(O"7604"), 16)), --             8#2035# => std_logic_vector(resize(unsigned'(O"0061"), 16)), --             8#2036# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2037# => std_logic_vector(resize(unsigned'(O"1061"), 16)), --             8#2040# => std_logic_vector(resize(unsigned'(O"7040"), 16)), --             8#2041# => std_logic_vector(resize(unsigned'(O"7450"), 16)), --             8#2042# => std_logic_vector(resize(unsigned'(O"5615"), 16)), --             8#2043# => std_logic_vector(resize(unsigned'(O"5614"), 16)), --             8#2044# => std_logic_vector(resize(unsigned'(O"2020"), 16)), --             8#2045# => std_logic_vector(resize(unsigned'(O"2001"), 16)), --             8#2046# => std_logic_vector(resize(unsigned'(O"2000"), 16)), --             8#2047# => std_logic_vector(resize(unsigned'(O"2074"), 16)), --             8#2050# => std_logic_vector(resize(unsigned'(O"2200"), 16)), --             8#2051# => std_logic_vector(resize(unsigned'(O"2075"), 16)), --             8#2052# => std_logic_vector(resize(unsigned'(O"2464"), 16)), --             8#2053# => std_logic_vector(resize(unsigned'(O"2465"), 16)), --             8#2054# => std_logic_vector(resize(unsigned'(O"2650"), 16)), --             8#2055# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2056# => std_logic_vector(resize(unsigned'(O"4026"), 16)), --             8#2057# => std_logic_vector(resize(unsigned'(O"4714"), 16)), --             8#2060# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2061# => std_logic_vector(resize(unsigned'(O"1056"), 16)), --             8#2062# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#2063# => std_logic_vector(resize(unsigned'(O"5266"), 16)), --             8#2064# => std_logic_vector(resize(unsigned'(O"4715"), 16)), --             8#2065# => std_logic_vector(resize(unsigned'(O"5655"), 16)), --             8#2066# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2067# => std_logic_vector(resize(unsigned'(O"1254"), 16)), --             8#2070# => std_logic_vector(resize(unsigned'(O"3714"), 16)), --             8#2071# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#2072# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2073# => std_logic_vector(resize(unsigned'(O"1075"), 16)), --             8#2074# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2075# => std_logic_vector(resize(unsigned'(O"1076"), 16)), --             8#2076# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2077# => std_logic_vector(resize(unsigned'(O"1077"), 16)), --             8#2100# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2101# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#2102# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2103# => std_logic_vector(resize(unsigned'(O"1053"), 16)), --             8#2104# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#2105# => std_logic_vector(resize(unsigned'(O"5716"), 16)), --             8#2106# => std_logic_vector(resize(unsigned'(O"4717"), 16)), --             8#2107# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#2110# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#2111# => std_logic_vector(resize(unsigned'(O"1052"), 16)), --             8#2112# => std_logic_vector(resize(unsigned'(O"3057"), 16)), --             8#2113# => std_logic_vector(resize(unsigned'(O"5720"), 16)), --             8#2114# => std_logic_vector(resize(unsigned'(O"2600"), 16)), --             8#2115# => std_logic_vector(resize(unsigned'(O"2732"), 16)), --             8#2116# => std_logic_vector(resize(unsigned'(O"2676"), 16)), --             8#2117# => std_logic_vector(resize(unsigned'(O"2702"), 16)), --             8#2120# => std_logic_vector(resize(unsigned'(O"2616"), 16)), --             8#2121# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2122# => std_logic_vector(resize(unsigned'(O"1245"), 16)), --             8#2123# => std_logic_vector(resize(unsigned'(O"3214"), 16)), --             8#2124# => std_logic_vector(resize(unsigned'(O"5234"), 16)), --             8#2125# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#2126# => std_logic_vector(resize(unsigned'(O"1251"), 16)), --             8#2127# => std_logic_vector(resize(unsigned'(O"3214"), 16)), --             8#2130# => std_logic_vector(resize(unsigned'(O"5234"), 16)), --             8#3000# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3001# => std_logic_vector(resize(unsigned'(O"1101"), 16)), --             8#3002# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3003# => std_logic_vector(resize(unsigned'(O"1076"), 16)), --             8#3004# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3005# => std_logic_vector(resize(unsigned'(O"1100"), 16)), --             8#3006# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3007# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#3010# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3011# => std_logic_vector(resize(unsigned'(O"4361"), 16)), --             8#3012# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#3013# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3014# => std_logic_vector(resize(unsigned'(O"1051"), 16)), --             8#3015# => std_logic_vector(resize(unsigned'(O"3057"), 16)), --             8#3016# => std_logic_vector(resize(unsigned'(O"4231"), 16)), --             8#3017# => std_logic_vector(resize(unsigned'(O"0137"), 16)), --             8#3020# => std_logic_vector(resize(unsigned'(O"3112"), 16)), --             8#3021# => std_logic_vector(resize(unsigned'(O"2112"), 16)), --             8#3022# => std_logic_vector(resize(unsigned'(O"7410"), 16)), --             8#3023# => std_logic_vector(resize(unsigned'(O"5600"), 16)), --             8#3024# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3025# => std_logic_vector(resize(unsigned'(O"1057"), 16)), --             8#3026# => std_logic_vector(resize(unsigned'(O"0410"), 16)), --             8#3027# => std_logic_vector(resize(unsigned'(O"4237"), 16)), --             8#3030# => std_logic_vector(resize(unsigned'(O"5221"), 16)), --             8#3031# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3032# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3033# => std_logic_vector(resize(unsigned'(O"1074"), 16)), --             8#3034# => std_logic_vector(resize(unsigned'(O"3010"), 16)), --             8#3035# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3036# => std_logic_vector(resize(unsigned'(O"5631"), 16)), --             8#3037# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3040# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#3041# => std_logic_vector(resize(unsigned'(O"5244"), 16)), --             8#3042# => std_logic_vector(resize(unsigned'(O"4302"), 16)), --             8#3043# => std_logic_vector(resize(unsigned'(O"5637"), 16)), --             8#3044# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3045# => std_logic_vector(resize(unsigned'(O"0106"), 16)), --             8#3046# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3047# => std_logic_vector(resize(unsigned'(O"5637"), 16)), --             8#3050# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3051# => std_logic_vector(resize(unsigned'(O"1273"), 16)), --             8#3052# => std_logic_vector(resize(unsigned'(O"3200"), 16)), --             8#3053# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#3054# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3055# => std_logic_vector(resize(unsigned'(O"1075"), 16)), --             8#3056# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3057# => std_logic_vector(resize(unsigned'(O"1076"), 16)), --             8#3060# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3061# => std_logic_vector(resize(unsigned'(O"4323"), 16)), --             8#3062# => std_logic_vector(resize(unsigned'(O"1055"), 16)), --             8#3063# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#3064# => std_logic_vector(resize(unsigned'(O"5307"), 16)), --             8#3065# => std_logic_vector(resize(unsigned'(O"4302"), 16)), --             8#3066# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#3067# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3070# => std_logic_vector(resize(unsigned'(O"1054"), 16)), --             8#3071# => std_logic_vector(resize(unsigned'(O"3057"), 16)), --             8#3072# => std_logic_vector(resize(unsigned'(O"5216"), 16)), --             8#3073# => std_logic_vector(resize(unsigned'(O"2465"), 16)), --             8#3074# => std_logic_vector(resize(unsigned'(O"2507"), 16)), --             8#3075# => std_logic_vector(resize(unsigned'(O"2744"), 16)), --             8#3076# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3077# => std_logic_vector(resize(unsigned'(O"0106"), 16)), --             8#3100# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3101# => std_logic_vector(resize(unsigned'(O"5674"), 16)), --             8#3102# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3103# => std_logic_vector(resize(unsigned'(O"7240"), 16)), --             8#3104# => std_logic_vector(resize(unsigned'(O"0105"), 16)), --             8#3105# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3106# => std_logic_vector(resize(unsigned'(O"5702"), 16)), --             8#3107# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3110# => std_logic_vector(resize(unsigned'(O"1106"), 16)), --             8#3111# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3112# => std_logic_vector(resize(unsigned'(O"5266"), 16)), --             8#3113# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3114# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3115# => std_logic_vector(resize(unsigned'(O"4041"), 16)), --             8#3116# => std_logic_vector(resize(unsigned'(O"1075"), 16)), --             8#3117# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3120# => std_logic_vector(resize(unsigned'(O"1100"), 16)), --             8#3121# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3122# => std_logic_vector(resize(unsigned'(O"5713"), 16)), --             8#3123# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3124# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3125# => std_logic_vector(resize(unsigned'(O"1075"), 16)), --             8#3126# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3127# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#3130# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3131# => std_logic_vector(resize(unsigned'(O"5723"), 16)), --             8#3132# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3133# => std_logic_vector(resize(unsigned'(O"1275"), 16)), --             8#3134# => std_logic_vector(resize(unsigned'(O"3200"), 16)), --             8#3135# => std_logic_vector(resize(unsigned'(O"4313"), 16)), --             8#3136# => std_logic_vector(resize(unsigned'(O"4323"), 16)), --             8#3137# => std_logic_vector(resize(unsigned'(O"1055"), 16)), --             8#3140# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#3141# => std_logic_vector(resize(unsigned'(O"5307"), 16)), --             8#3142# => std_logic_vector(resize(unsigned'(O"4302"), 16)), --             8#3143# => std_logic_vector(resize(unsigned'(O"5266"), 16)), --             8#3144# => std_logic_vector(resize(unsigned'(O"7200"), 16)), --             8#3145# => std_logic_vector(resize(unsigned'(O"1273"), 16)), --             8#3146# => std_logic_vector(resize(unsigned'(O"3200"), 16)), --             8#3147# => std_logic_vector(resize(unsigned'(O"4313"), 16)), --             8#3150# => std_logic_vector(resize(unsigned'(O"1077"), 16)), --             8#3151# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3152# => std_logic_vector(resize(unsigned'(O"1102"), 16)), --             8#3153# => std_logic_vector(resize(unsigned'(O"4020"), 16)), --             8#3154# => std_logic_vector(resize(unsigned'(O"1053"), 16)), --             8#3155# => std_logic_vector(resize(unsigned'(O"7440"), 16)), --             8#3156# => std_logic_vector(resize(unsigned'(O"5276"), 16)), --             8#3157# => std_logic_vector(resize(unsigned'(O"4302"), 16)), --             8#3160# => std_logic_vector(resize(unsigned'(O"5674"), 16)), --             8#3161# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3162# => std_logic_vector(resize(unsigned'(O"1140"), 16)), --             8#3163# => std_logic_vector(resize(unsigned'(O"4237"), 16)), --             8#3164# => std_logic_vector(resize(unsigned'(O"5761"), 16)), --             8#3165# => std_logic_vector(resize(unsigned'(O"2146"), 16)), --             8#0200# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0201# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0202# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0203# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0204# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0205# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0206# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0207# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0210# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0211# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0212# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0213# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0214# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0215# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0216# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0217# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0220# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0221# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0222# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0223# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0224# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0225# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0226# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0227# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0230# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0231# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0232# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0233# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0234# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0235# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0236# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0237# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0240# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0241# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0242# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0243# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0244# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0245# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0246# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0247# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0250# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0251# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0252# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0253# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0254# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#0255# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3400# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3401# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3402# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3403# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3404# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3405# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3406# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3407# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3410# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3411# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3412# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3413# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3414# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3415# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3416# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3417# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3420# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3421# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3422# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3423# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3424# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3425# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3426# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3427# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3430# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3431# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3432# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3433# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3434# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3435# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3436# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3437# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3440# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3441# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3442# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3443# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3444# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3445# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3446# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3447# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3450# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3451# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3452# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3453# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3454# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3455# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3456# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3457# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3460# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3461# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3462# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3463# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3464# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3465# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3466# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3467# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3470# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3471# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3472# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3473# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3474# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3475# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3476# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#3477# => std_logic_vector(resize(unsigned'(O"0252"), 16)), --             8#2652# => std_logic_vector(resize(unsigned'(O"3203"), 16)), --             8#2653# => std_logic_vector(resize(unsigned'(O"3371"), 16)), --             8#2654# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2655# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2656# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2657# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2660# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2661# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2662# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2663# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2664# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2665# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2666# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2667# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2670# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2671# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2672# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2673# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2674# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2675# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2676# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2677# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2700# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2701# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2702# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2703# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2704# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2705# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2706# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2707# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2710# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2711# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2712# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2713# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2714# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2715# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2716# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2717# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2720# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2721# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2722# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2723# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2724# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2725# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2726# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2727# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2730# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2731# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2732# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2733# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2734# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2735# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2736# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2737# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2740# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2741# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2742# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             8#2743# => std_logic_vector(resize(unsigned'(O"0000"), 16)), --             others  => X"0000"
       );
	attribute syn_ramstyle : string;
	attribute syn_ramstyle of ramdata : signal is "block_ram";
    signal raddr : integer range 0 to 4095 := 0;
begin
    Q <= ramdata(raddr);

    process (Clock, Reset) is
    begin
        if Reset = '1' then
            raddr <= 0;
        elsif rising_edge(Clock) then
            if ClockEn = '1' then 
                raddr <= to_integer(unsigned(Address));
                if WE = '1' then 
                    ramdata(to_integer(unsigned(Address))) <= Data;
                end if;
            end if;
        end if;
    end process;

end architecture logic;

